* Two Stage Single Slope ADC using skywater 130nm

.lib "models/sky130.lib.spice" ff
.lib adc_sky.lib nops_noprot

xadc_a vref vin clock reset vdd gnd xout yout ADC_ANALOG
* comparator xout rises with clock when it does rise. and falls with it too
* comparator yout does the same but is inverted in terms of the comparison
* both should be read on falling edge

* Input Signals

Vdd vdd GND 1.8
V5  clock GND PULSE(0 1.8 0 10p 10p .5u 1u)
Vin vin GND 0.5
V2  GND vref 1
V3  reset GND PULSE(0 1.8 0 10p 10p 20n 256.02u)


.option method=Gear
.ic v(xadc_a.inp)=0

.control
set color0=white

let vdelta = 1/256
let dstart = 0
let dstop  = 256
let num_sim= 256

let vstart = dstart * vdelta
let vstop  = dstop * vdelta
let ddelta = (dstop - dstart)/num_sim
*let vdelta = (vstop-vstart)/num_sim
let vact   = vstart
let dact   = dstart

set ext = "v.txt"
set dlm = "_"

shell mkdir -p outfiles/sky
set wr_singlescale
set wr_vecnames

while vact < vstop
    echo
    echo Running Sweep $&dact/$&dstop
    echo
    alter vin vact
    ;run
    tran 1u 512u uic

    let cut-tstart = 256u
    let cut-tstop = 512u
    cutout

    ;plot I(vdd)
    wrdata outfiles/sky_raw_d$&dact$ext -I(vdd)

    let lin-tstart = 256u
    let lin-tstop  = 512u
    let lin-tstep  = 100n
    linearize I(vdd)

    ;plot I(vdd)
    wrdata outfiles/sky_lin_d$&dact$ext -I(vdd)

    let dact = dact + ddelta
    let vact = dact * vdelta

    destroy all
end
*exit
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
