* Two Stage Single Slope ADC using skywater 130nm

.lib "models/sky130.lib.spice" $corner
.lib "adc_sky.lib"             nops_noprot ;$flavor
.inc "adc_wrap.cir"

xadc vin vref clock reset vdda vddd gnd d7 d6 d5 d4 d3 d2 d1 d0 ADC_WRAP 
        
Vdda vdda   GND   1.8
Vddd vddd   GND   1.8
V5   clock  GND   PULSE(0 1.8 0 10p 10p .5u 1u)
Vin  vin    GND   0.5
V2   GND    vref  1
V3   reset  GND   PULSE(0 1.8 0 10p 10p 20n 256.02u)

.option method=Gear
.ic v(xadc.xanalog.inp)=0

.control
set color0=white

let vdelta = 1/256
let dstart = $start
let dstop  = $stop
let num_sim= $count

let vstart = dstart * vdelta
let vstop  = dstop * vdelta
let ddelta = (dstop - dstart)/num_sim
*let vdelta = (vstop-vstart)/num_sim
let vact   = vstart
let dact   = dstart

set ext = "v.txt"
set dlm = "_"

${iswrite}shell mkdir -p ../outfiles/sky
set wr_singlescale
set wr_vecnames
    
while vact < vstop
    echo
    echo Running Sweep $&dact/$&dstop
    echo
    alter vin vact
    ;run
    tran 1u 512u uic

    let cut-tstart = 256u
    let cut-tstop = 512u
    cutout

    ${isplot} plot I(vdd)
    ${iswrite}wrdata outfiles/sky_raw_d$&dact$ext -I(vddd) -I(vdda)

    let lin-tstart = 256u
    let lin-tstop  = 512u
    let lin-tstep  = 100n
    linearize I(vdd)

    ${isplot} plot I(vdd)
    ${iswrite}wrdata outfiles/sky_lin_d$&dact$ext -I(vddd) -I(vdda)

    let dact = dact + ddelta
    let vact = dact * vdelta

    ${isbatch}destroy all
end
${isbatch}exit
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
