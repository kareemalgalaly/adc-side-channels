* Single slope adc
*.include lib/lmx58_lm2904.lib
.include adc.lib

* Parameters

.param vdd=3.3
.param vss=0
.param per={1u}
.param rise={per/5}

* Supplies / References

vdd   vdd   gnd {vdd}
vin   vin   gnd  1
vref  vref  gnd -1

* Control Signals

vclk     clock   gnd PULSE({vss} {vdd} {per/2}  {rise} {rise} {per/2} {per})
vrestart restart gnd PULSE({vss} {vdd} {per*10} {rise} {rise} {per}   {per*256})
vresetn  resetn  gnd PWL(0 {vss}, {per*8}, {vss}, {per*8.2}, {vdd})

* DUT

*xcore vin vref comp_out restart resetn vdd gnd ADC_CORE r=250 c={330n}
xadc vin vref clock resetn restart d7 d6 d5 d4 d3 d2 d1 d0 vdd gnd ADC vdd={vdd} vss={vss}

r7 d7 gnd 1k
r6 d6 gnd 1k
r5 d5 gnd 1k
r4 d4 gnd 1k
r3 d3 gnd 1k
r2 d2 gnd 1k
r1 d1 gnd 1k
r0 d0 gnd 1k

.options TRTOL=1.0 CHGTOL=1e-16 ; switches near caps

.control
*tran 10n 550u uic
*tran 100n 550u

* adc_core
* plot V(vin) V(comp_out) V(xcore.ramp_out) V(restart)
* plot V(resetn) V(restart)

;plot V(vin) V(xadc.comp_out) V(xadc.xcore.ramp_out) V(restart)
;plot -I(vdd)
let vstart = 1
let vstop  = 3.3
let vdelta = 4.0
let vact   = vstart

while vact <= vstop
    echo Running Sweep $&vact/$&vstop
    echo
    alter vin vact
    ;run
    tran 10n 550u uic

    let digitized=(V(d0) + V(d1)*2 + V(d2)*4 + V(d3)*8 + V(d4)*16 + V(d5)*32 + V(d6)*64 + V(d7))*128
    ;plot digitized -I(vdd)

    linearize I(vdd) digitized

    meas tran teval WHEN digitized=0.001 RISE=1
    echo Start point $&teval
    let cut-tstart = teval

    meas tran teval WHEN digitized=0.001 FALL=1
    echo End point $&teval
    let cut-tstop = teval

    cutout


    plot I(vdd) digitized

    set wr_singlescale
    set wr_vecnames
    wrdata out.txt -I(vdd) digitized
    set appendwrite

    let vact = vact + vdelta
end

;plot tran1.digitized tran2.digitized tran3.digitized
plot I(tran1.vdd) I(tran2.vdd) I(tran3.vdd)
.endc

.end
