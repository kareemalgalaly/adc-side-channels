* Two Stage Single Slope ADC using skywater 130nm

.lib "models/sky130.lib.spice" tt
.lib adc_sky.lib nops_noprot

xadc_a vref vin clock reset vdd gnd xout yout ADC_ANALOG
* comparator xout rises with clock when it does rise. and falls with it too
* comparator yout does the same but is inverted in terms of the comparison
* both should be read on falling edge

* Input Signals

Vdd vdd GND 1.8
V5  clock GND PULSE(0 1.8 0 10p 10p .5u 1u)
Vin vin GND 0.5
V2  GND vref 1
V3  reset GND PULSE(0 1.8 0 10p 10p 20n 256.02u)


.option method=Gear
.ic v(xadc_a.inp)=0

.control
set color0=white

let vstart = 0
let vstop  = 1.0
let num_sim= 1
let vdelta = (vstop-vstart)/num_sim
let vact   = vstart
let digit  = 0

set ext = "v.txt"
set dlm = "_"

while vact < vstop
    echo
    echo Running Sweep $&digit/$&num_sim
    echo
    alter vin vact
    ;run
    tran 1u 512u uic

    let lin-tstart = 257u
    let lin-tstop  = 512u
    let lin-tstep  = 100n

    plot I(vdd)
    ; linearize I(vdd) ; digitized
    ; plot I(vdd)

    let cut-tstart = 257u
    let cut-tstop = 512u
    cutout

    set wr_singlescale
    set wr_vecnames
    wrdata ../outfiles/sky/sky_d$&digit$dlm$&vact$ext -I(vdd) ;digitized

    let vact = vact + vdelta
    let digit = digit + 1

    ;destroy all
end
*exit
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
