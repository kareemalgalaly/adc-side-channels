* Single slope adc
*.include lib/lmx58_lm2904.lib
*.include ~/Documents/SpiceLibraries/LT/ADI_ng.lib
*.include ~/Documents/SpiceLibraries/kareem.lib
.include adc.lib

* Parameters

.param vdd=3.3
.param vss=0
.param per={1u}
.param rise={per/10}

* Supplies / References

vdd   vdd   gnd {vdd}
vin   vin   gnd  1
vref  vref  gnd -1

* Control Signals

vclk     clock   gnd PULSE({vss} {vdd} {per/2}  {rise} {rise} {per/2} {per})
vrestart restart gnd PULSE({vss} {vdd} {per*10} {rise} {rise} {per}   {per*256})
vresetn  resetn  gnd PWL(0 {vss}, {per*8}, {vss}, {per*8.2}, {vdd})

* DUT

*xadc vin vref resetn restart 7 6 5 4 3 2 1 0 vdd vss ADC vdd={vdd} vss={vss}
xcore vin vref comp_out restart resetn vdd gnd ADC_CORE r=250 c={330n}

.options TRTOL=1.0 CHGTOL=1e-16 ; switches near caps

.control
tran 10n 550u uic
*tran 100n 550u

* adc_core
plot V(vin) V(comp_out) V(xcore.ramp_out) V(restart)
plot V(resetn) V(restart)

*let digitized=(V(0)/128 + V(1)/64 + V(2)/32 + V(3)/16 + V(4)/8 + V(5)/4 + V(6)/2 + V(7))/13.2+0.5
*plot digitized
*plot V(vin) V(xadc.xcore.ramp_out) V(xadc.comp_out)
plot -I(vdd)



*linearize I(vdd)
*wrdata out.txt I(vdd)
.endc

.end
