* Two Stage Single Slope ADC using skywater 130nm

.lib "models/sky130.lib.spice" $corner
.lib "adc_sky.lib"             nops_noprot ;$flavor
.inc "adc_wrap.cir"

xadc vin vref clock reset vdda vddd gnd d7 d6 d5 d4 d3 d2 d1 d0 ADC_WRAP 
        
Vdda vdda   GND   1.8
Vddd vddd   GND   1.8
V5   clock  GND   PULSE(0 1.8 0 10p 10p .5u 1u)
Vin  vin    GND   0.5
V2   GND    vref  1
V3   reset  GND   PULSE(0 1.8 0 10p 10p 20n 256.02u)

.option method=Gear
.ic v(xadc.xanalog.inp)=0

.control
set color0=white

let vstart = $vstart
let vstop  = $vstop
let num_sim= $vcount
let vdelta = (vstop-vstart)/num_sim
let vact   = vstart
let digit  = 0

set ext = "v.txt"
set dlm = "_"

while vact < vstop
    echo
    echo Running Sweep $&digit/$&num_sim
    echo
    alter vin vact
    ;run
    tran 1u 512u uic

    let lin-tstart = 257u
    let lin-tstop  = 512u
    let lin-tstep  = 100n

    ${isplot}${islin} plot -I(vdda) -I(vddd)
    ${islin}          linearize I(vdda) I(vddd) ; digitized
    ${isplot}         plot -I(vdda) -I(vddd)

    let cut-tstart = 257u
    let cut-tstop = 512u
    cutout
    ;plot -I(vdda) -I(vddd)

    set wr_singlescale
    set wr_vecnames
    ${iswrite}wrdata ../outfiles/sky/sky_d$&digit$dlm$&vact$ext -I(vddd) -I(vdda) ;digitized

    let vact = vact + vdelta
    let digit = digit + 1

    ${isbatch}destroy all
end
${isbatch}exit
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
