* NMOS Transfer and Output Characteristics
* Generated 10-Oct-2021 10:31:26
* Include SkyWater sky130 device models

.lib "models/sky130.lib.spice" tt

.option scale=1e-6

xm1 d1 g1 0 0   sky130_fd_pr__nfet_01v8_lvt w=1 l=0.5
vgs g1 0        dc=0.9
vds d1 0        dc=0.9

.control
dc vgs 0 1.8 0.01
*wrdata nmos_01v8_transfer_tt.dat -i(vds)
plot title "VGS" -i(vds)

dc vds 0 1.8 0.01
*wrdata nmos_01v8_output_tt.dat -i(vds)
plot title "VDS" -i(vds)
.endc

.end

