* Single slope adc
.include ../lib/adc.lib

* Parameters

.param vdd=3.3
.param vss=0
.param per={1u}
.param rise={per/5}

* Supplies / References

vdd   vdd   gnd {vdd}
rdd   vdd   gnd 1e6
vin   vin   gnd  1
rin   vin   gnd 1e6
vref  vref  gnd -1
rref  vref  gnd 1e6

* Control Signals

vclk     clock   gnd PULSE({vss} {vdd} {per/2}  {rise} {rise} {per/2} {per})
vrestart restart gnd PULSE({vss} {vdd} {per*10} {rise} {rise} {per}   {per*256})
vresetn  resetn  gnd PWL(0 {vss}, {per*8}, {vss}, {per*8.2}, {vdd})

* DUT

*xcore vin vref comp_out restart resetn vdd gnd ADC_CORE r=250 c={330n}
xadc vin vref clock resetn restart d7 d6 d5 d4 d3 d2 d1 d0 vdd gnd ADC vdd={vdd} vss={vss}

r7 d7 gnd 1k
r6 d6 gnd 1k
r5 d5 gnd 1k
r4 d4 gnd 1k
r3 d3 gnd 1k
r2 d2 gnd 1k
r1 d1 gnd 1k
r0 d0 gnd 1k

.options TRTOL=1.0 CHGTOL=1e-16 ; switches near caps

.control

let vstart = 0
let vstop  = 3.3
let vdelta = 1.0
let vact   = vstart

while vact <= vstop
    echo Running Sweep $&vact/$&vstop
    echo
    alter vin vact
    ;run
    tran 10n 550u uic

    let digitized=(V(d0) + V(d1)*2 + V(d2)*4 + V(d3)*8 + V(d4)*16 + V(d5)*32 + V(d6)*64 + V(d7))*128

    plot -I(vdd) digitized*2e-7 ; V(restart)*2m
    linearize I(vdd) digitized V(restart)

    let cut-tstart = 10u
    let cut-tstop = 266u

    cutout

    set wr_singlescale
    set wr_vecnames
    wrdata ../outfiles/out_$&vact -I(vdd) digitized
    set appendwrite

    let vact = vact + vdelta
end
.endc

.end
