* Single slope adc using comp w/ preamp
.lib "models/sky130.lib.spice" tt
.include ../lib/adc.lib
.include ../lib/comp_ceyda.spice

.param vdd=1.8
.param vss=0
.param vmid={vdd/2}
.param per={1u}
.param rise={per/5}

* Supplies / References

vdd   vdd   gnd {vdd}
rdd   vdd   gnd 1e6
vin   vin   gnd  1
rin   vin   gnd 1e6
vref  vref  gnd -1
rref  vref  gnd 1e6

* Control Signals

vclk     clock   gnd PULSE({vss} {vdd} {per/2}  {rise} {rise} {per/2} {per})
vrestart restart gnd PULSE({vss} {vdd} {per*10} {rise} {rise} {per}   {per*256})
vresetn  resetn  gnd PWL(0 {vss}, {per*8}, {vss}, {per*8.2}, {vdd})


xramp vref vramp reset enable vdd gnd RAMP_GEN r=100 c=1u
xcomp vramp vin   clock  vdd gnd comp_outp comp_outn COMP

* Digital Components
a_dig_ctrl [d_clk d_resetn d_comp_out d_start_over] [d_ramp_reset d_enable d_busy d_valid d7 d6 d5 d4 d3 d2 d1 d0] null dmodel
.model dmodel d_cosim simulation="../../build/adc.so"

* Interface
abridge_a [clock resetn comp_outp restart] [d_clk d_resetn d_comp_out d_start_over] auto_adc
abridge_d [d_ramp_reset d_enable d_busy d_valid d7 d6 d5 d4 d3 d2 d1 d0] [rreset enable busy valid v7 v6 v5 v4 v3 v2 v1 v0] auto_dac
.model auto_adc adc_bridge(in_low  = {vdd/2}    in_high  = {vdd/2})
*.model auto_adc adc_bridge(in_low  = {vdd/2-.1}  in_high  = {vdd/2+.1})
.model auto_dac dac_bridge(out_low = 0          out_high = {vdd})

.control
tran 10n 550u uic
plot V(vin) V(vdd) V(vramp) V(comp_outp)
.endc

.end
