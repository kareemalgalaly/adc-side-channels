* NGSPICE file created from latch_2_pex.ext - technology: sky130A

.subckt latch_2 vdd ck out1 out2 in2 in1 vss
X0 a_1257_3075.t8 ck.t0 vdd.t17 vdd.t16 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_698_3956.t11 in2.t0 a_2200_588.t9 vss.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=9e+06u l=900000u
X2 a_1257_3075.t4 a_1315_3049.t15 a_772_588.t11 vss.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=9e+06u l=900000u
X3 a_2200_588.t8 in2.t1 a_698_3956.t10 vss.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=9e+06u l=900000u
X4 a_1257_3075.t11 a_1315_3049.t16 vdd.t31 vdd.t30 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=900000u
X5 vdd.t5 a_1257_3075.t15 a_1315_3049.t14 vdd.t4 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=900000u
X6 a_1257_3075.t12 a_1315_3049.t17 vdd.t33 vdd.t32 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=900000u
X7 vdd.t1 a_1315_3049.t18 a_1257_3075.t0 vdd.t0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=900000u
X8 a_1257_3075.t1 a_1315_3049.t19 a_772_588.t10 vss.t1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=9e+06u l=900000u
X9 out2.t1 a_1315_3049.t20 vdd.t29 vdd.t28 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 vdd.t21 a_1257_3075.t16 a_1315_3049.t13 vdd.t20 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=900000u
X11 a_1315_3049.t8 a_1257_3075.t17 a_2200_588.t17 vss.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=9e+06u l=900000u
X12 a_1315_3049.t12 a_1257_3075.t18 vdd.t23 vdd.t22 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=900000u
X13 a_1315_3049.t11 a_1257_3075.t19 vdd.t25 vdd.t24 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=900000u
X14 vdd.t15 ck.t1 a_1315_3049.t0 vdd.t14 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_1315_3049.t7 a_1257_3075.t20 a_2200_588.t12 vss.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=9e+06u l=900000u
X16 a_772_588.t9 a_1315_3049.t21 a_1257_3075.t9 vss.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=9e+06u l=900000u
X17 a_698_3956.t9 in2.t2 a_2200_588.t5 vss.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=9e+06u l=900000u
X18 out2.t0 a_1315_3049.t22 vss.t6 vss.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X19 a_2200_588.t4 in2.t3 a_698_3956.t8 vss.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=9e+06u l=900000u
X20 a_1315_3049.t10 a_1257_3075.t21 vdd.t19 vdd.t18 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=900000u
X21 vdd.t9 a_1257_3075.t22 out1.t1 vdd.t8 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_698_3956.t7 in2.t4 a_2200_588.t1 vss.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=9e+06u l=900000u
X23 a_698_3956.t15 in1.t0 a_772_588.t13 vss.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=9e+06u l=900000u
X24 a_2200_588.t0 in2.t5 a_698_3956.t6 vss.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=9e+06u l=900000u
X25 a_698_3956.t5 in2.t6 a_2200_588.t3 vss.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=9e+06u l=900000u
X26 vdd.t13 ck.t2 a_772_588.t2 vdd.t12 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_772_588.t8 a_1315_3049.t23 a_1257_3075.t5 vss.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=9e+06u l=900000u
X28 a_2200_588.t11 a_1257_3075.t23 a_1315_3049.t6 vss.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=9e+06u l=900000u
X29 a_698_3956.t4 in2.t7 a_2200_588.t2 vss.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=9e+06u l=900000u
X30 a_1257_3075.t2 a_1315_3049.t24 vdd.t3 vdd.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=900000u
X31 vss.t20 ck.t3 a_698_3956.t12 vss.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=900000u
X32 a_1315_3049.t5 a_1257_3075.t24 a_2200_588.t14 vss.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=9e+06u l=900000u
X33 a_772_588.t3 in1.t1 a_698_3956.t13 vss.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=9e+06u l=900000u
X34 a_1257_3075.t3 a_1315_3049.t25 a_772_588.t7 vss.t2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=9e+06u l=900000u
X35 a_2200_588.t13 a_1257_3075.t25 a_1315_3049.t4 vss.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=9e+06u l=900000u
X36 vdd.t35 a_1315_3049.t26 a_1257_3075.t13 vdd.t34 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=900000u
X37 a_1257_3075.t14 a_1315_3049.t27 a_772_588.t6 vss.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=9e+06u l=900000u
X38 a_1315_3049.t3 a_1257_3075.t26 a_2200_588.t16 vss.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=9e+06u l=900000u
X39 a_2200_588.t7 in2.t8 a_698_3956.t3 vss.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=9e+06u l=900000u
X40 vdd.t27 a_1257_3075.t27 a_1315_3049.t9 vdd.t26 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=900000u
X41 a_772_588.t14 in1.t2 a_698_3956.t16 vss.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=9e+06u l=900000u
X42 a_2200_588.t10 ck.t4 vdd.t11 vdd.t10 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X43 vss.t30 a_1257_3075.t28 out1.t0 vss.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X44 a_698_3956.t18 in1.t3 a_772_588.t16 vss.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=9e+06u l=900000u
X45 a_772_588.t5 a_1315_3049.t28 a_1257_3075.t6 vss.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=9e+06u l=900000u
X46 a_2200_588.t15 a_1257_3075.t29 a_1315_3049.t2 vss.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=9e+06u l=900000u
X47 a_698_3956.t17 in1.t4 a_772_588.t15 vss.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=9e+06u l=900000u
X48 a_772_588.t18 in1.t5 a_698_3956.t20 vss.t41 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=9e+06u l=900000u
X49 a_698_3956.t19 in1.t6 a_772_588.t17 vss.t40 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=9e+06u l=900000u
X50 a_772_588.t12 in1.t7 a_698_3956.t14 vss.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=9e+06u l=900000u
X51 a_698_3956.t0 in1.t8 a_772_588.t0 vss.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=9e+06u l=900000u
X52 a_772_588.t1 in1.t9 a_698_3956.t1 vss.t3 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=9e+06u l=900000u
X53 vdd.t7 a_1315_3049.t29 a_1257_3075.t7 vdd.t6 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=900000u
X54 a_2200_588.t6 in2.t9 a_698_3956.t2 vss.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=9e+06u l=900000u
X55 a_772_588.t4 a_1315_3049.t30 a_1257_3075.t10 vss.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=9e+06u l=900000u
X56 a_2200_588.t18 a_1257_3075.t30 a_1315_3049.t1 vss.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=9e+06u l=900000u
R0 ck.t4 ck.t1 558.241
R1 ck.t0 ck.t2 552.833
R2 ck.n1 ck.t4 248.438
R3 ck.n0 ck.t0 245.261
R4 ck.n0 ck.t3 124.659
R5 ck.n1 ck.n0 3.35
R6 ck ck.n1 0.002
R7 vdd.n71 vdd.n70 347.481
R8 vdd.n148 vdd.n145 272.304
R9 vdd.n137 vdd.n136 234.277
R10 vdd.n78 vdd.n77 226.529
R11 vdd.n119 vdd.n111 201.018
R12 vdd.n138 vdd.n137 185.574
R13 vdd.n115 vdd.n114 185
R14 vdd.n101 vdd.n100 185
R15 vdd.n91 vdd.n90 185
R16 vdd.n77 vdd.n76 185
R17 vdd.n1 vdd.n0 185
R18 vdd.n23 vdd.n18 172.799
R19 vdd.t6 vdd.t2 144.196
R20 vdd.t32 vdd.t6 144.196
R21 vdd.t26 vdd.t18 144.196
R22 vdd.t24 vdd.t4 144.196
R23 vdd.t34 vdd.t30 144.196
R24 vdd.n101 vdd.n99 143.811
R25 vdd.n24 vdd.n23 132.893
R26 vdd.n52 vdd.n51 121.599
R27 vdd.n116 vdd.n115 115.952
R28 vdd.n109 vdd.n108 115.199
R29 vdd.n7 vdd.n6 108.046
R30 vdd.n3 vdd.t20 90.88
R31 vdd.n134 vdd.n133 84.215
R32 vdd.t2 vdd.n2 81.792
R33 vdd.n42 vdd.n39 79.811
R34 vdd.n106 vdd.t16 71.473
R35 vdd.n21 vdd.t28 71.473
R36 vdd.n21 vdd.t8 71.473
R37 vdd.n96 vdd.t12 68.495
R38 vdd.n140 vdd.n92 66.039
R39 vdd.t12 vdd.n95 64.345
R40 vdd.n44 vdd.t10 64.028
R41 vdd.n146 vdd.t24 58.769
R42 vdd.n134 vdd.t0 47.863
R43 vdd.n4 vdd.t14 40.203
R44 vdd.n143 vdd.t34 39.987
R45 vdd.n142 vdd.n91 36.369
R46 vdd.n102 vdd.t17 32.505
R47 vdd.n102 vdd.t13 32.505
R48 vdd.n30 vdd.t29 32.505
R49 vdd.n30 vdd.t9 32.505
R50 vdd.n43 vdd.t11 32.505
R51 vdd.n43 vdd.t15 32.505
R52 vdd.n103 vdd.n101 28.009
R53 vdd.n46 vdd.n42 26.823
R54 vdd.n54 vdd.n9 23.824
R55 vdd.n74 vdd.n73 23.628
R56 vdd.n78 vdd.n1 22.4
R57 vdd.n74 vdd.t32 15.146
R58 vdd.n73 vdd.n3 14.54
R59 vdd.n137 vdd.t22 13.934
R60 vdd.n125 vdd.n124 13.176
R61 vdd.n94 vdd.n93 9.3
R62 vdd.n78 vdd.n75 9.3
R63 vdd.n75 vdd.n74 9.3
R64 vdd.n133 vdd.n132 9.088
R65 vdd.n59 vdd.n58 8.854
R66 vdd.n105 vdd.n97 7.058
R67 vdd.n92 vdd.t26 6.058
R68 vdd.n82 vdd.t3 4.76
R69 vdd.n82 vdd.t7 4.76
R70 vdd.n83 vdd.t33 4.76
R71 vdd.n83 vdd.t21 4.76
R72 vdd.n85 vdd.t19 4.76
R73 vdd.n85 vdd.t27 4.76
R74 vdd.n80 vdd.t23 4.76
R75 vdd.n80 vdd.t35 4.76
R76 vdd.n79 vdd.t31 4.76
R77 vdd.n79 vdd.t1 4.76
R78 vdd.n88 vdd.t25 4.76
R79 vdd.n88 vdd.t5 4.76
R80 vdd.n148 vdd.n142 4.616
R81 vdd.n123 vdd.n122 4.094
R82 vdd.n60 vdd.n59 4.093
R83 vdd.n32 vdd.n31 3.148
R84 vdd.n106 vdd.n96 2.978
R85 vdd.n84 vdd.n82 1.695
R86 vdd.n81 vdd.n79 1.645
R87 vdd.n47 vdd.n46 1.6
R88 vdd.n54 vdd.n10 1.489
R89 vdd.n39 vdd.n38 1.217
R90 vdd.n38 vdd.n37 1.217
R91 vdd.n132 vdd.n94 1.211
R92 vdd.n84 vdd.n83 1.206
R93 vdd.n86 vdd.n85 1.195
R94 vdd.n81 vdd.n80 1.189
R95 vdd.n89 vdd.n88 1.166
R96 vdd.n149 vdd.n78 1.069
R97 vdd vdd.n89 0.897
R98 vdd.n103 vdd.n102 0.786
R99 vdd.n104 vdd.n103 0.731
R100 vdd.n46 vdd.n43 0.704
R101 vdd.n87 vdd.n86 0.515
R102 vdd.n87 vdd.n81 0.51
R103 vdd.n86 vdd.n84 0.51
R104 vdd.n31 vdd.n30 0.452
R105 vdd vdd.n149 0.443
R106 vdd.n124 vdd.n123 0.29
R107 vdd.n120 vdd.n110 0.244
R108 vdd.n110 vdd.n109 0.244
R109 vdd.n126 vdd.n125 0.244
R110 vdd.n132 vdd.n126 0.244
R111 vdd.n149 vdd.n148 0.225
R112 vdd.n148 vdd 0.187
R113 vdd.n59 vdd.n57 0.134
R114 vdd.n42 vdd.n41 0.127
R115 vdd.n41 vdd.n40 0.127
R116 vdd.n53 vdd.n52 0.125
R117 vdd.n54 vdd.n53 0.125
R118 vdd.n6 vdd.n5 0.109
R119 vdd.n5 vdd.n4 0.109
R120 vdd.n135 vdd.n134 0.073
R121 vdd.n136 vdd.n135 0.067
R122 vdd.n25 vdd.n24 0.066
R123 vdd.n26 vdd.n25 0.066
R124 vdd.n16 vdd.n15 0.064
R125 vdd.n26 vdd.n16 0.064
R126 vdd.n69 vdd.n68 0.06
R127 vdd.n70 vdd.n69 0.06
R128 vdd.n55 vdd.n8 0.058
R129 vdd.n8 vdd.n7 0.058
R130 vdd.n118 vdd.n117 0.045
R131 vdd.n117 vdd.n116 0.045
R132 vdd.n36 vdd.n35 0.039
R133 vdd.n37 vdd.n36 0.039
R134 vdd.n48 vdd.n47 0.037
R135 vdd.n49 vdd.n48 0.037
R136 vdd.n106 vdd.n105 0.037
R137 vdd.n105 vdd.n104 0.037
R138 vdd.n28 vdd.n27 0.035
R139 vdd.n29 vdd.n28 0.035
R140 vdd.n46 vdd.n45 0.028
R141 vdd.n45 vdd.n44 0.028
R142 vdd.n34 vdd.n12 0.025
R143 vdd.n56 vdd.n55 0.025
R144 vdd.n118 vdd.n113 0.025
R145 vdd.n27 vdd.n14 0.025
R146 vdd.n113 vdd.n112 0.025
R147 vdd.n14 vdd.n13 0.025
R148 vdd.n12 vdd.n11 0.025
R149 vdd.n57 vdd.n56 0.025
R150 vdd.n108 vdd.n107 0.019
R151 vdd.n107 vdd.n106 0.019
R152 vdd.n23 vdd.n22 0.019
R153 vdd.n22 vdd.n21 0.019
R154 vdd.n20 vdd.n19 0.019
R155 vdd.n21 vdd.n20 0.019
R156 vdd.n51 vdd.n50 0.019
R157 vdd.n50 vdd.n49 0.019
R158 vdd.n99 vdd.n98 0.013
R159 vdd.n18 vdd.n17 0.013
R160 vdd.n34 vdd.n33 0.009
R161 vdd.n33 vdd.n32 0.009
R162 vdd.n66 vdd.n63 0.008
R163 vdd.n121 vdd.n120 0.008
R164 vdd.n122 vdd.n121 0.008
R165 vdd.n63 vdd.n62 0.008
R166 vdd.n131 vdd.n130 0.007
R167 vdd.n68 vdd.n61 0.007
R168 vdd.n130 vdd.n129 0.007
R169 vdd.n61 vdd.n60 0.007
R170 vdd.n66 vdd.n65 0.006
R171 vdd.n131 vdd.n128 0.006
R172 vdd.n128 vdd.n127 0.006
R173 vdd.n72 vdd.n71 0.006
R174 vdd.n73 vdd.n72 0.006
R175 vdd.n145 vdd.n144 0.006
R176 vdd.n144 vdd.n143 0.006
R177 vdd.n65 vdd.n64 0.006
R178 vdd.n148 vdd.n147 0.006
R179 vdd.n147 vdd.n146 0.006
R180 vdd.n139 vdd.n138 0.002
R181 vdd.n140 vdd.n139 0.002
R182 vdd.n142 vdd.n141 0.002
R183 vdd.n141 vdd.n140 0.002
R184 vdd.n31 vdd.n29 0.001
R185 vdd.n27 vdd.n26 0.001
R186 vdd.n120 vdd.n119 0.001
R187 vdd.n55 vdd.n54 0.001
R188 vdd.n119 vdd.n118 0.001
R189 vdd.n89 vdd.n87 0.001
R190 vdd.n68 vdd.n67 0.001
R191 vdd.n37 vdd.n34 0.001
R192 vdd.n132 vdd.n131 0.001
R193 vdd.n67 vdd.n66 0.001
R194 a_1257_3075.n15 a_1257_3075.t17 312.468
R195 a_1257_3075.n21 a_1257_3075.t30 255.73
R196 a_1257_3075.n20 a_1257_3075.t24 255.73
R197 a_1257_3075.n19 a_1257_3075.t23 255.73
R198 a_1257_3075.n18 a_1257_3075.t20 255.73
R199 a_1257_3075.n17 a_1257_3075.t29 255.73
R200 a_1257_3075.n16 a_1257_3075.t26 255.73
R201 a_1257_3075.n15 a_1257_3075.t25 255.73
R202 a_1257_3075.n8 a_1257_3075.t22 244.213
R203 a_1257_3075.n3 a_1257_3075.t16 240.005
R204 a_1257_3075.n0 a_1257_3075.t18 239.261
R205 a_1257_3075.n5 a_1257_3075.t19 177.833
R206 a_1257_3075.n4 a_1257_3075.t27 177.833
R207 a_1257_3075.n3 a_1257_3075.t21 177.833
R208 a_1257_3075.n0 a_1257_3075.t15 160.666
R209 a_1257_3075.n8 a_1257_3075.t28 152.018
R210 a_1257_3075.n4 a_1257_3075.n3 62.171
R211 a_1257_3075.n5 a_1257_3075.n4 62.171
R212 a_1257_3075.n16 a_1257_3075.n15 56.738
R213 a_1257_3075.n17 a_1257_3075.n16 56.738
R214 a_1257_3075.n18 a_1257_3075.n17 56.738
R215 a_1257_3075.n19 a_1257_3075.n18 56.738
R216 a_1257_3075.n20 a_1257_3075.n19 56.738
R217 a_1257_3075.n21 a_1257_3075.n20 56.738
R218 a_1257_3075.n6 a_1257_3075.n5 55.787
R219 a_1257_3075.n13 a_1257_3075.t8 33.499
R220 a_1257_3075.n9 a_1257_3075.n8 6.998
R221 a_1257_3075.n14 a_1257_3075.n13 5.775
R222 a_1257_3075.n7 a_1257_3075.n0 5.547
R223 a_1257_3075.n9 a_1257_3075.t2 4.761
R224 a_1257_3075.n12 a_1257_3075.t0 4.761
R225 a_1257_3075.n2 a_1257_3075.t13 4.76
R226 a_1257_3075.n2 a_1257_3075.t11 4.76
R227 a_1257_3075.n10 a_1257_3075.t7 4.76
R228 a_1257_3075.n10 a_1257_3075.t12 4.76
R229 a_1257_3075.n22 a_1257_3075.n21 4.033
R230 a_1257_3075.n1 a_1257_3075.n7 3.865
R231 a_1257_3075.n14 a_1257_3075.t9 3.147
R232 a_1257_3075.n1 a_1257_3075.n11 2.688
R233 a_1257_3075.n22 a_1257_3075.t14 1.934
R234 a_1257_3075.n23 a_1257_3075.t6 1.933
R235 a_1257_3075.n23 a_1257_3075.t4 1.933
R236 a_1257_3075.n25 a_1257_3075.t5 1.933
R237 a_1257_3075.n25 a_1257_3075.t3 1.933
R238 a_1257_3075.n28 a_1257_3075.t10 1.933
R239 a_1257_3075.t1 a_1257_3075.n28 1.933
R240 a_1257_3075.n24 a_1257_3075.n22 1.508
R241 a_1257_3075.n26 a_1257_3075.n25 1.217
R242 a_1257_3075.n28 a_1257_3075.n27 1.208
R243 a_1257_3075.n11 a_1257_3075.n9 1.161
R244 a_1257_3075.n24 a_1257_3075.n23 1.156
R245 a_1257_3075.n12 a_1257_3075.n1 1.153
R246 a_1257_3075.n13 a_1257_3075.n12 0.885
R247 a_1257_3075.n1 a_1257_3075.n2 0.657
R248 a_1257_3075.n11 a_1257_3075.n10 0.65
R249 a_1257_3075.n7 a_1257_3075.n6 0.453
R250 a_1257_3075.n27 a_1257_3075.n14 0.31
R251 a_1257_3075.n26 a_1257_3075.n24 0.308
R252 a_1257_3075.n27 a_1257_3075.n26 0.303
R253 in2.n4 in2.t9 337.009
R254 in2.n0 in2.t7 331.236
R255 in2.n7 in2.t3 255.758
R256 in2.n6 in2.t2 255.758
R257 in2.n5 in2.t1 255.758
R258 in2.n4 in2.t0 255.758
R259 in2.n3 in2.t4 255.758
R260 in2.n2 in2.t5 255.758
R261 in2.n1 in2.t6 255.758
R262 in2.n0 in2.t8 255.758
R263 in2.n7 in2.n6 82.044
R264 in2.n5 in2.n4 81.252
R265 in2.n6 in2.n5 81.252
R266 in2.n1 in2.n0 75.478
R267 in2.n2 in2.n1 75.478
R268 in2.n3 in2.n2 75.478
R269 in2.n8 in2.n3 42.505
R270 in2.n8 in2.n7 41.369
R271 in2 in2.n8 0.568
R272 a_2200_588.n0 a_2200_588.t10 36.414
R273 a_2200_588.n12 a_2200_588.t2 1.933
R274 a_2200_588.n12 a_2200_588.t7 1.933
R275 a_2200_588.n4 a_2200_588.t1 1.933
R276 a_2200_588.n4 a_2200_588.t4 1.933
R277 a_2200_588.n2 a_2200_588.t5 1.933
R278 a_2200_588.n2 a_2200_588.t8 1.933
R279 a_2200_588.n1 a_2200_588.t9 1.933
R280 a_2200_588.n1 a_2200_588.t6 1.933
R281 a_2200_588.n7 a_2200_588.t16 1.933
R282 a_2200_588.n7 a_2200_588.t15 1.933
R283 a_2200_588.n6 a_2200_588.t12 1.933
R284 a_2200_588.n6 a_2200_588.t11 1.933
R285 a_2200_588.n10 a_2200_588.t14 1.933
R286 a_2200_588.n10 a_2200_588.t18 1.933
R287 a_2200_588.n0 a_2200_588.t17 1.933
R288 a_2200_588.n0 a_2200_588.t13 1.933
R289 a_2200_588.n15 a_2200_588.t3 1.933
R290 a_2200_588.t0 a_2200_588.n15 1.933
R291 a_2200_588.n13 a_2200_588.n11 1.54
R292 a_2200_588.n3 a_2200_588.n1 1.238
R293 a_2200_588.n8 a_2200_588.n0 1.166
R294 a_2200_588.n13 a_2200_588.n12 1.145
R295 a_2200_588.n3 a_2200_588.n2 0.917
R296 a_2200_588.n15 a_2200_588.n14 0.909
R297 a_2200_588.n5 a_2200_588.n4 0.893
R298 a_2200_588.n11 a_2200_588.n10 0.732
R299 a_2200_588.n9 a_2200_588.n6 0.73
R300 a_2200_588.n8 a_2200_588.n7 0.727
R301 a_2200_588.n11 a_2200_588.n9 0.414
R302 a_2200_588.n9 a_2200_588.n8 0.399
R303 a_2200_588.n5 a_2200_588.n3 0.374
R304 a_2200_588.n14 a_2200_588.n5 0.372
R305 a_2200_588.n14 a_2200_588.n13 0.099
R306 a_698_3956.n0 a_698_3956.t12 11.545
R307 a_698_3956.n14 a_698_3956.t8 1.933
R308 a_698_3956.n14 a_698_3956.t9 1.933
R309 a_698_3956.n12 a_698_3956.t6 1.933
R310 a_698_3956.n12 a_698_3956.t7 1.933
R311 a_698_3956.n6 a_698_3956.t1 1.933
R312 a_698_3956.n6 a_698_3956.t19 1.933
R313 a_698_3956.n8 a_698_3956.t16 1.933
R314 a_698_3956.n8 a_698_3956.t4 1.933
R315 a_698_3956.n10 a_698_3956.t3 1.933
R316 a_698_3956.n10 a_698_3956.t5 1.933
R317 a_698_3956.n5 a_698_3956.t20 1.933
R318 a_698_3956.n5 a_698_3956.t18 1.933
R319 a_698_3956.n2 a_698_3956.t14 1.933
R320 a_698_3956.n2 a_698_3956.t17 1.933
R321 a_698_3956.n1 a_698_3956.t2 1.933
R322 a_698_3956.n1 a_698_3956.t0 1.933
R323 a_698_3956.n0 a_698_3956.t13 1.933
R324 a_698_3956.n0 a_698_3956.t15 1.933
R325 a_698_3956.n17 a_698_3956.t10 1.933
R326 a_698_3956.t11 a_698_3956.n17 1.933
R327 a_698_3956.n7 a_698_3956.n6 1.899
R328 a_698_3956.n3 a_698_3956.n0 1.869
R329 a_698_3956.n17 a_698_3956.n16 1.474
R330 a_698_3956.n3 a_698_3956.n2 1.457
R331 a_698_3956.n13 a_698_3956.n12 1.455
R332 a_698_3956.n4 a_698_3956.n1 1.454
R333 a_698_3956.n11 a_698_3956.n10 1.446
R334 a_698_3956.n7 a_698_3956.n5 1.437
R335 a_698_3956.n15 a_698_3956.n14 1.423
R336 a_698_3956.n9 a_698_3956.n8 1.423
R337 a_698_3956.n9 a_698_3956.n7 0.405
R338 a_698_3956.n11 a_698_3956.n9 0.401
R339 a_698_3956.n16 a_698_3956.n15 0.4
R340 a_698_3956.n13 a_698_3956.n11 0.398
R341 a_698_3956.n16 a_698_3956.n4 0.396
R342 a_698_3956.n4 a_698_3956.n3 0.392
R343 a_698_3956.n15 a_698_3956.n13 0.358
R344 vss.n79 vss.n77 20291
R345 vss.n85 vss.n74 20088.2
R346 vss.n89 vss.n78 13987
R347 vss.n92 vss.n91 13784.2
R348 vss.n86 vss.n83 1305.22
R349 vss.n93 vss.n72 888.341
R350 vss.n88 vss.n87 835.173
R351 vss.n87 vss.n78 585
R352 vss.n67 vss.n66 585
R353 vss.n84 vss.n78 522.992
R354 vss.t40 vss.t3 485.264
R355 vss.t41 vss.t40 485.264
R356 vss.t38 vss.t41 485.264
R357 vss.t24 vss.t38 485.264
R358 vss.t10 vss.t24 485.264
R359 vss.t9 vss.t10 485.264
R360 vss.t11 vss.t9 485.264
R361 vss.t12 vss.t11 485.264
R362 vss.t13 vss.t12 485.264
R363 vss.t15 vss.t14 485.264
R364 vss.t16 vss.t15 485.264
R365 vss.t17 vss.t16 485.264
R366 vss.t8 vss.t17 485.264
R367 vss.t0 vss.t8 485.264
R368 vss.t22 vss.t0 485.264
R369 vss.t37 vss.t22 485.264
R370 vss.t21 vss.t37 485.264
R371 vss.t23 vss.t21 485.264
R372 vss.t4 vss.t18 485.264
R373 vss.t7 vss.t4 485.264
R374 vss.t2 vss.t26 485.264
R375 vss.t26 vss.t1 485.264
R376 vss.t36 vss.t32 485.264
R377 vss.t28 vss.t31 485.264
R378 vss.t35 vss.t34 485.264
R379 vss.t34 vss.t33 485.264
R380 vss.n9 vss.t39 475.076
R381 vss.n15 vss.t25 475.069
R382 vss.n3 vss.n2 438.907
R383 vss.n81 vss.n80 418.347
R384 vss.n37 vss.n10 417.81
R385 vss.n87 vss.n86 409.975
R386 vss.n80 vss.n71 407.636
R387 vss.n59 vss.t5 406.153
R388 vss.n59 vss.t29 406.153
R389 vss.n0 vss.t27 327.361
R390 vss.n84 vss.t23 325.476
R391 vss.n41 vss.t36 311.955
R392 vss.n38 vss.n3 286.216
R393 vss.n22 vss.n17 279.34
R394 vss.n27 vss.n15 260.049
R395 vss.n35 vss.t7 242.632
R396 vss.n35 vss.t2 242.632
R397 vss.n6 vss.t28 242.632
R398 vss.t3 vss.n73 240.594
R399 vss.n75 vss.t13 240.593
R400 vss.n38 vss.t35 240.593
R401 vss.n79 vss.n73 226.334
R402 vss.n91 vss.n74 208.588
R403 vss.t14 vss.n76 169.23
R404 vss.n23 vss.n22 165.646
R405 vss.n47 vss.n41 163.113
R406 vss.n61 vss.n56 150.587
R407 vss.n85 vss.n84 145.83
R408 vss.n1 vss.n0 144.036
R409 vss.n62 vss.n61 73.479
R410 vss.n90 vss.n76 73.401
R411 vss.n63 vss.n53 69.487
R412 vss.n54 vss.t6 39.6
R413 vss.n54 vss.t30 39.6
R414 vss.n68 vss.n67 23.532
R415 vss.n83 vss.n72 13.552
R416 vss.n82 vss.n77 9.3
R417 vss.n77 vss.n75 9.3
R418 vss.n95 vss.n94 9.3
R419 vss.n71 vss.n69 9.3
R420 vss.n81 vss.n70 7.899
R421 vss.n36 vss.n31 6.277
R422 vss.n94 vss.n71 5.894
R423 vss.n89 vss.n77 5.794
R424 vss.n31 vss.t20 4.892
R425 vss.n82 vss.n81 4.19
R426 vss.n38 vss.n37 2.537
R427 vss.n37 vss.n36 2.101
R428 vss.n90 vss.n75 2.038
R429 vss.n65 vss.n38 1.928
R430 vss.n62 vss.n54 1.781
R431 vss.n65 vss.n64 1.13
R432 vss.n94 vss.n93 0.673
R433 vss vss.n68 0.397
R434 vss vss.n95 0.348
R435 vss.n88 vss.n82 0.345
R436 vss.n38 vss.n8 0.317
R437 vss.n31 vss.n30 0.26
R438 vss.n64 vss.n63 0.127
R439 vss.n24 vss.n23 0.105
R440 vss.n27 vss.n24 0.105
R441 vss.n26 vss.n25 0.104
R442 vss.n27 vss.n26 0.104
R443 vss.n64 vss.n50 0.065
R444 vss.n56 vss.n55 0.061
R445 vss.n53 vss.n52 0.061
R446 vss.n52 vss.n51 0.061
R447 vss.n61 vss.n60 0.059
R448 vss.n60 vss.n59 0.059
R449 vss.n59 vss.n58 0.059
R450 vss.n58 vss.n57 0.059
R451 vss.n48 vss.n40 0.055
R452 vss.n40 vss.n39 0.055
R453 vss.n49 vss.n48 0.053
R454 vss.n50 vss.n49 0.053
R455 vss.n19 vss.n18 0.049
R456 vss.t19 vss.n19 0.049
R457 vss.n22 vss.n21 0.049
R458 vss.n21 vss.n20 0.041
R459 vss.n28 vss.n12 0.031
R460 vss.n95 vss.n69 0.031
R461 vss.n12 vss.n11 0.031
R462 vss.n46 vss.n45 0.02
R463 vss.n45 vss.n44 0.02
R464 vss.n17 vss.n16 0.016
R465 vss.n46 vss.n43 0.014
R466 vss.n43 vss.n42 0.014
R467 vss.n63 vss.n62 0.013
R468 vss.n7 vss.n6 0.013
R469 vss.n8 vss.n7 0.013
R470 vss.n92 vss.n73 0.011
R471 vss.n93 vss.n69 0.011
R472 vss.n93 vss.n92 0.011
R473 vss.n20 vss.t19 0.009
R474 vss.n14 vss.n13 0.007
R475 vss.n86 vss.n85 0.007
R476 vss.n80 vss.n79 0.007
R477 vss.n15 vss.n14 0.007
R478 vss.n10 vss.n9 0.007
R479 vss.n2 vss.n1 0.007
R480 vss.n33 vss.n32 0.007
R481 vss.n5 vss.n4 0.007
R482 vss.n6 vss.n5 0.007
R483 vss.n83 vss.n74 0.005
R484 vss.n76 vss.n74 0.005
R485 vss.n91 vss.n72 0.005
R486 vss.n91 vss.n90 0.005
R487 vss.n90 vss.n89 0.005
R488 vss.n89 vss.n88 0.005
R489 vss.n34 vss.n33 0.004
R490 vss.n35 vss.n34 0.004
R491 vss.n94 vss.n70 0.002
R492 vss.n29 vss.n28 0.001
R493 vss.n70 vss.n69 0.001
R494 vss.n30 vss.n29 0.001
R495 vss.n68 vss.n65 0.001
R496 vss.n28 vss.n27 0.001
R497 vss.n48 vss.n47 0.001
R498 vss.n47 vss.n46 0.001
R499 vss.n36 vss.n35 0.001
R500 a_1315_3049.n13 a_1315_3049.t21 317.901
R501 a_1315_3049.n19 a_1315_3049.t27 255.73
R502 a_1315_3049.n18 a_1315_3049.t28 255.73
R503 a_1315_3049.n17 a_1315_3049.t15 255.73
R504 a_1315_3049.n16 a_1315_3049.t23 255.73
R505 a_1315_3049.n15 a_1315_3049.t25 255.73
R506 a_1315_3049.n14 a_1315_3049.t30 255.73
R507 a_1315_3049.n13 a_1315_3049.t19 255.73
R508 a_1315_3049.n10 a_1315_3049.t20 243.336
R509 a_1315_3049.n8 a_1315_3049.t24 240.005
R510 a_1315_3049.n3 a_1315_3049.t18 239.064
R511 a_1315_3049.n3 a_1315_3049.t16 177.833
R512 a_1315_3049.n8 a_1315_3049.t29 177.833
R513 a_1315_3049.n9 a_1315_3049.t17 168.114
R514 a_1315_3049.n4 a_1315_3049.t26 160.713
R515 a_1315_3049.n10 a_1315_3049.t22 152.811
R516 a_1315_3049.n19 a_1315_3049.n18 62.171
R517 a_1315_3049.n18 a_1315_3049.n17 62.171
R518 a_1315_3049.n17 a_1315_3049.n16 62.171
R519 a_1315_3049.n16 a_1315_3049.n15 62.171
R520 a_1315_3049.n15 a_1315_3049.n14 62.171
R521 a_1315_3049.n14 a_1315_3049.n13 62.171
R522 a_1315_3049.n4 a_1315_3049.n3 60.554
R523 a_1315_3049.n9 a_1315_3049.n8 50.114
R524 a_1315_3049.n11 a_1315_3049.t0 33.805
R525 a_1315_3049.n11 a_1315_3049.n10 5.168
R526 a_1315_3049.n6 a_1315_3049.t9 4.76
R527 a_1315_3049.n6 a_1315_3049.t11 4.76
R528 a_1315_3049.n2 a_1315_3049.t14 4.76
R529 a_1315_3049.n2 a_1315_3049.t12 4.76
R530 a_1315_3049.n1 a_1315_3049.t13 4.76
R531 a_1315_3049.n1 a_1315_3049.t10 4.76
R532 a_1315_3049.n5 a_1315_3049.n4 4.691
R533 a_1315_3049.t8 a_1315_3049.n27 3.296
R534 a_1315_3049.n12 a_1315_3049.n11 3.151
R535 a_1315_3049.n21 a_1315_3049.t1 2.949
R536 a_1315_3049.n21 a_1315_3049.n20 2.311
R537 a_1315_3049.n0 a_1315_3049.n9 2.054
R538 a_1315_3049.n22 a_1315_3049.t6 1.933
R539 a_1315_3049.n22 a_1315_3049.t5 1.933
R540 a_1315_3049.n24 a_1315_3049.t2 1.933
R541 a_1315_3049.n24 a_1315_3049.t7 1.933
R542 a_1315_3049.n26 a_1315_3049.t4 1.933
R543 a_1315_3049.n26 a_1315_3049.t3 1.933
R544 a_1315_3049.n12 a_1315_3049.n1 1.876
R545 a_1315_3049.n20 a_1315_3049.n12 1.772
R546 a_1315_3049.n25 a_1315_3049.n24 1.056
R547 a_1315_3049.n23 a_1315_3049.n22 1.023
R548 a_1315_3049.n27 a_1315_3049.n26 1.022
R549 a_1315_3049.n20 a_1315_3049.n19 0.736
R550 a_1315_3049.n5 a_1315_3049.n2 0.637
R551 a_1315_3049.n1 a_1315_3049.n0 0.616
R552 a_1315_3049.n7 a_1315_3049.n6 0.612
R553 a_1315_3049.n7 a_1315_3049.n5 0.558
R554 a_1315_3049.n0 a_1315_3049.n7 0.556
R555 a_1315_3049.n25 a_1315_3049.n23 0.309
R556 a_1315_3049.n27 a_1315_3049.n25 0.307
R557 a_1315_3049.n23 a_1315_3049.n21 0.292
R558 a_772_588.n0 a_772_588.t2 36.546
R559 a_772_588.n10 a_772_588.t13 3.235
R560 a_772_588.n4 a_772_588.t1 3.234
R561 a_772_588.n8 a_772_588.n6 2.938
R562 a_772_588.n2 a_772_588.t7 1.933
R563 a_772_588.n2 a_772_588.t4 1.933
R564 a_772_588.n1 a_772_588.t6 1.933
R565 a_772_588.n1 a_772_588.t5 1.933
R566 a_772_588.n0 a_772_588.t10 1.933
R567 a_772_588.n0 a_772_588.t9 1.933
R568 a_772_588.n9 a_772_588.t15 1.933
R569 a_772_588.n9 a_772_588.t3 1.933
R570 a_772_588.n5 a_772_588.t16 1.933
R571 a_772_588.n5 a_772_588.t14 1.933
R572 a_772_588.n3 a_772_588.t17 1.933
R573 a_772_588.n3 a_772_588.t18 1.933
R574 a_772_588.n7 a_772_588.t0 1.933
R575 a_772_588.n7 a_772_588.t12 1.933
R576 a_772_588.t11 a_772_588.n15 1.933
R577 a_772_588.n15 a_772_588.t8 1.933
R578 a_772_588.n12 a_772_588.n11 1.545
R579 a_772_588.n6 a_772_588.n5 0.939
R580 a_772_588.n8 a_772_588.n7 0.906
R581 a_772_588.n10 a_772_588.n9 0.905
R582 a_772_588.n4 a_772_588.n3 0.879
R583 a_772_588.n14 a_772_588.n1 0.868
R584 a_772_588.n13 a_772_588.n2 0.56
R585 a_772_588.n12 a_772_588.n0 0.533
R586 a_772_588.n15 a_772_588.n14 0.516
R587 a_772_588.n6 a_772_588.n4 0.388
R588 a_772_588.n14 a_772_588.n13 0.3
R589 a_772_588.n13 a_772_588.n12 0.287
R590 a_772_588.n11 a_772_588.n10 0.226
R591 a_772_588.n11 a_772_588.n8 0.154
R592 out2 out2.t0 40.768
R593 out2 out2.t1 33.755
R594 out1 out1.t0 40.556
R595 out1 out1.t1 33.768
R596 in1.n0 in1.t0 335.456
R597 in1.n4 in1.t9 331.809
R598 in1.n2 in1.t7 255.758
R599 in1.n1 in1.t4 255.758
R600 in1.n0 in1.t1 255.758
R601 in1.n6 in1.t3 255.758
R602 in1.n5 in1.t5 255.758
R603 in1.n4 in1.t6 255.758
R604 in1.n7 in1.t2 241.027
R605 in1.n3 in1.t8 241.022
R606 in1.n1 in1.n0 79.698
R607 in1.n2 in1.n1 79.698
R608 in1.n3 in1.n2 77.861
R609 in1.n5 in1.n4 75.478
R610 in1.n6 in1.n5 75.478
R611 in1.n7 in1.n6 74.181
R612 in1 in1.n7 19.506
R613 in1 in1.n3 16.996
C0 out1 out2 0.23fF
C1 vdd out1 0.83fF
C2 vdd out2 0.66fF
C3 in2 in1 0.36fF
C4 ck vdd 2.43fF
.ends

